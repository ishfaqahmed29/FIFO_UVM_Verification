import uvm_pkg::*;
`include "uvm_macros.svh"

// ----COVERAGE----

class fifo_coverage extends uvm_subscriber #(data_item);

    
        
    function new();
        
    endfunction: new 

endclass: fifo_coverage